* C:\Users\shesh\Desktop\DIGITAL CIRCUITS LABORATORY ASSIGNMENT\GRAY_TO_BINARY_CONVERTERS_USING_NAND_GATE\GRAY_TO_BINARY_CONVERTERS_USING_NAND_GATE.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 22 23:05:39 2020



** Analysis setup **
.tran 1ms 6ms
.OP 
.STMLIB "C:\Users\shesh\Documents\graytobinary.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "GRAY_TO_BINARY_CONVERTERS_USING_NAND_GATE.net"
.INC "GRAY_TO_BINARY_CONVERTERS_USING_NAND_GATE.als"


.probe


.END
