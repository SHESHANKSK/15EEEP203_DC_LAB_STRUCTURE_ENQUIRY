* C:\Users\shesh\Desktop\DIGITAL CIRCUITS LABORATORY ASSIGNMENT\HALF_SUBSTRACTOR_USING_74153_MULTIPLEXER\HALF_SUBSTRACTOR_USING_74153_MULTIPLEXER.sch

* Schematics Version 9.1 - Web Update 1
* Mon Nov 23 11:36:19 2020



** Analysis setup **
.tran 10ms 100ms
.OP 
.STMLIB "C:\Users\shesh\Desktop\DIGITAL CIRCUITS LABORATORY ASSIGNMENT\HALF_SUBSTRACTOR_USING_74153_MULTIPLEXER.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "HALF_SUBSTRACTOR_USING_74153_MULTIPLEXER.net"
.INC "HALF_SUBSTRACTOR_USING_74153_MULTIPLEXER.als"


.probe


.END
